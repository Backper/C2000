module dma_ctrl (
    input clk;
    input rstn;
);

reg [4:0]ps;
reg [4:0]ns;

always@(*)begin
    ns = IDLE;
    
end
    
endmodule